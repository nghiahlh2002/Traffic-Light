library verilog;
use verilog.vl_types.all;
entity traffic_tb is
end traffic_tb;
