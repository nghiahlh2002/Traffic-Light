library verilog;
use verilog.vl_types.all;
entity \time__vlg_vec_tst\ is
end \time__vlg_vec_tst\;
