library verilog;
use verilog.vl_types.all;
entity ngovao_vlg_vec_tst is
end ngovao_vlg_vec_tst;
